For this project we ae not using Full adder and ripple carry adder as a two dseperate verilog file 
   we are using only 1 verliog that is PES_RCA.v file which is there in the repo


// module PES_FA(A, B, clk, S, Cout);
	// input A, B, clk;
	// output S, Cout;

	// assign S = A ^ B;
	// assign Cout = A | B;
// endmodule
