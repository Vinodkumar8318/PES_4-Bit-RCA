For this project we ae not using Full adder and ripple carry adder as a 2 Seperate verilog files. 
  So We are using only 1 verliog and 1 Test bench file that is PES_RCA.v and PES_RCA_TB.v files which is there in the repo.


// module PES_FA(A, B, clk, S, Cout);
	// input A, B, clk;
	// output S, Cout;

	// assign S = A ^ B;
	// assign Cout = A | B;
// endmodule
